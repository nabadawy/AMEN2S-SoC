module iota (
	input in_st_0,
	input rndc_r,
	output out_st_0
);

assign out_st_0 = in_st_0 ^ rndc_r;


endmodule
